module testbench (
	input         clock,
	input         reset,

	output        io_dmem_invalidate_lr,
	input         io_dmem_ordered,
	input         io_dmem_replay_next,
	output [39:0] io_dmem_req_bits_addr,
	output [4:0]  io_dmem_req_bits_cmd,
	output        io_dmem_req_bits_phys,
	output [6:0]  io_dmem_req_bits_tag,
	output [2:0]  io_dmem_req_bits_typ,
	input         io_dmem_req_ready,
	output        io_dmem_req_valid,
	input  [63:0] io_dmem_resp_bits_data,
	input  [63:0] io_dmem_resp_bits_data_word_bypass,
	input         io_dmem_resp_bits_has_data,
	input         io_dmem_resp_bits_replay,
	input  [6:0]  io_dmem_resp_bits_tag,
	input  [2:0]  io_dmem_resp_bits_typ,
	input         io_dmem_resp_valid,
	output [63:0] io_dmem_s1_data_data,
	output [7:0]  io_dmem_s1_data_mask,
	output        io_dmem_s1_kill,
	input         io_dmem_s2_nack,
	input         io_dmem_s2_xcpt_ae_ld,
	input         io_dmem_s2_xcpt_ae_st,
	input         io_dmem_s2_xcpt_ma_ld,
	input         io_dmem_s2_xcpt_ma_st,
	input         io_dmem_s2_xcpt_pf_ld,
	input         io_dmem_s2_xcpt_pf_st,

	input         io_fpu_dec_ren1,
	input         io_fpu_dec_ren2,
	input         io_fpu_dec_ren3,
	input         io_fpu_dec_wen,
	output [63:0] io_fpu_dmem_resp_data,
	output [4:0]  io_fpu_dmem_resp_tag,
	output [2:0]  io_fpu_dmem_resp_type,
	output        io_fpu_dmem_resp_val,
	input  [4:0]  io_fpu_fcsr_flags_bits,
	input         io_fpu_fcsr_flags_valid,
	input         io_fpu_fcsr_rdy,
	output [2:0]  io_fpu_fcsr_rm,
	output [63:0] io_fpu_fromint_data,
	input         io_fpu_illegal_rm,
	output [31:0] io_fpu_inst,
	output        io_fpu_killm,
	output        io_fpu_killx,
	input         io_fpu_nack_mem,
	input         io_fpu_sboard_clr,
	input  [4:0]  io_fpu_sboard_clra,
	input         io_fpu_sboard_set,
	input  [63:0] io_fpu_store_data,
	input  [63:0] io_fpu_toint_data,
	output        io_fpu_valid,

	input         io_hartid,

	output        io_imem_bht_update_bits_mispredict,
	output [38:0] io_imem_bht_update_bits_pc,
	output [6:0]  io_imem_bht_update_bits_prediction_bits_bht_history,
	output [1:0]  io_imem_bht_update_bits_prediction_bits_bht_value,
	output        io_imem_bht_update_bits_prediction_valid,
	output        io_imem_bht_update_bits_taken,
	output        io_imem_bht_update_valid,
	output [38:0] io_imem_btb_update_bits_br_pc,
	output [1:0]  io_imem_btb_update_bits_cfiType,
	output        io_imem_btb_update_bits_isValid,
	output [38:0] io_imem_btb_update_bits_pc,
	output [6:0]  io_imem_btb_update_bits_prediction_bits_bht_history,
	output [1:0]  io_imem_btb_update_bits_prediction_bits_bht_value,
	output [5:0]  io_imem_btb_update_bits_prediction_bits_entry,
	output        io_imem_btb_update_bits_prediction_valid,
	output        io_imem_btb_update_valid,
	output        io_imem_flush_icache,
	output [39:0] io_imem_req_bits_pc,
	output        io_imem_req_bits_speculative,
	output        io_imem_req_valid,
	input         io_imem_resp_bits_ae,
	input  [6:0]  io_imem_resp_bits_btb_bits_bht_history,
	input  [1:0]  io_imem_resp_bits_btb_bits_bht_value,
	input         io_imem_resp_bits_btb_bits_bridx,
	input  [5:0]  io_imem_resp_bits_btb_bits_entry,
	input         io_imem_resp_bits_btb_bits_taken,
	input         io_imem_resp_bits_btb_valid,
	input  [31:0] io_imem_resp_bits_data,
	input  [39:0] io_imem_resp_bits_pc,
	input         io_imem_resp_bits_pf,
	input         io_imem_resp_bits_replay,
	output        io_imem_resp_ready,
	input         io_imem_resp_valid,
	output        io_imem_sfence_bits_rs1,
	output        io_imem_sfence_bits_rs2,
	output        io_imem_sfence_valid,

	input         io_interrupts_debug,
	input         io_interrupts_meip,
	input         io_interrupts_msip,
	input         io_interrupts_mtip,
	input         io_interrupts_seip,

	output        io_ptw_invalidate,
	output [29:0] io_ptw_pmp_0_addr,
	output [1:0]  io_ptw_pmp_0_cfg_a,
	output        io_ptw_pmp_0_cfg_l,
	output        io_ptw_pmp_0_cfg_r,
	output        io_ptw_pmp_0_cfg_w,
	output        io_ptw_pmp_0_cfg_x,
	output [31:0] io_ptw_pmp_0_mask,
	output [29:0] io_ptw_pmp_1_addr,
	output [1:0]  io_ptw_pmp_1_cfg_a,
	output        io_ptw_pmp_1_cfg_l,
	output        io_ptw_pmp_1_cfg_r,
	output        io_ptw_pmp_1_cfg_w,
	output        io_ptw_pmp_1_cfg_x,
	output [31:0] io_ptw_pmp_1_mask,
	output [29:0] io_ptw_pmp_2_addr,
	output [1:0]  io_ptw_pmp_2_cfg_a,
	output        io_ptw_pmp_2_cfg_l,
	output        io_ptw_pmp_2_cfg_r,
	output        io_ptw_pmp_2_cfg_w,
	output        io_ptw_pmp_2_cfg_x,
	output [31:0] io_ptw_pmp_2_mask,
	output [29:0] io_ptw_pmp_3_addr,
	output [1:0]  io_ptw_pmp_3_cfg_a,
	output        io_ptw_pmp_3_cfg_l,
	output        io_ptw_pmp_3_cfg_r,
	output        io_ptw_pmp_3_cfg_w,
	output        io_ptw_pmp_3_cfg_x,
	output [31:0] io_ptw_pmp_3_mask,
	output [29:0] io_ptw_pmp_4_addr,
	output [1:0]  io_ptw_pmp_4_cfg_a,
	output        io_ptw_pmp_4_cfg_l,
	output        io_ptw_pmp_4_cfg_r,
	output        io_ptw_pmp_4_cfg_w,
	output        io_ptw_pmp_4_cfg_x,
	output [31:0] io_ptw_pmp_4_mask,
	output [29:0] io_ptw_pmp_5_addr,
	output [1:0]  io_ptw_pmp_5_cfg_a,
	output        io_ptw_pmp_5_cfg_l,
	output        io_ptw_pmp_5_cfg_r,
	output        io_ptw_pmp_5_cfg_w,
	output        io_ptw_pmp_5_cfg_x,
	output [31:0] io_ptw_pmp_5_mask,
	output [29:0] io_ptw_pmp_6_addr,
	output [1:0]  io_ptw_pmp_6_cfg_a,
	output        io_ptw_pmp_6_cfg_l,
	output        io_ptw_pmp_6_cfg_r,
	output        io_ptw_pmp_6_cfg_w,
	output        io_ptw_pmp_6_cfg_x,
	output [31:0] io_ptw_pmp_6_mask,
	output [29:0] io_ptw_pmp_7_addr,
	output [1:0]  io_ptw_pmp_7_cfg_a,
	output        io_ptw_pmp_7_cfg_l,
	output        io_ptw_pmp_7_cfg_r,
	output        io_ptw_pmp_7_cfg_w,
	output        io_ptw_pmp_7_cfg_x,
	output [31:0] io_ptw_pmp_7_mask,
	output [15:0] io_ptw_ptbr_asid,
	output [3:0]  io_ptw_ptbr_mode,
	output [43:0] io_ptw_ptbr_ppn,
	output [1:0]  io_ptw_status_dprv,
	output        io_ptw_status_mxr,
	output [1:0]  io_ptw_status_prv,
	output        io_ptw_status_sum,

	input         io_rocc_cmd_ready,
	output        io_rocc_cmd_valid,
	input         io_rocc_interrupt
);
	wire [31:0] rvfi_insn;
	wire [63:0] rvfi_mem_addr;
	wire [63:0] rvfi_mem_rdata;
	wire [7:0]  rvfi_mem_rmask;
	wire [63:0] rvfi_mem_wdata;
	wire [7:0]  rvfi_mem_wmask;
	wire [7:0]  rvfi_order;
	wire [63:0] rvfi_pc_rdata;
	wire [63:0] rvfi_pc_wdata;
	wire [4:0]  rvfi_rd_addr;
	wire [63:0] rvfi_rd_wdata;
	wire [4:0]  rvfi_rs1_addr;
	wire [63:0] rvfi_rs1_rdata;
	wire [4:0]  rvfi_rs2_addr;
	wire [63:0] rvfi_rs2_rdata;
	wire        rvfi_trap;
	wire        rvfi_valid;

	reg [7:0] insn_count = 0;
	reg [7:0] cycle_count = 0;

	always @(posedge clock) begin
		if (!reset && rvfi_valid)
			insn_count <= insn_count + |(insn_count + 1);
		cycle_count <= cycle_count + |(cycle_count + 1);
	end

	always @* begin
		assume(reset == (cycle_count < 5));
		cover(insn_count == 1);
		cover(insn_count == 2);
		cover(insn_count == 3);
		cover(insn_count == 4);
	end

	RocketWithRVFI uut (
		.clock                                              (clock                                              ),
		.io_dmem_invalidate_lr                              (io_dmem_invalidate_lr                              ),
		.io_dmem_ordered                                    (io_dmem_ordered                                    ),
		.io_dmem_replay_next                                (io_dmem_replay_next                                ),
		.io_dmem_req_bits_addr                              (io_dmem_req_bits_addr                              ),
		.io_dmem_req_bits_cmd                               (io_dmem_req_bits_cmd                               ),
		.io_dmem_req_bits_phys                              (io_dmem_req_bits_phys                              ),
		.io_dmem_req_bits_tag                               (io_dmem_req_bits_tag                               ),
		.io_dmem_req_bits_typ                               (io_dmem_req_bits_typ                               ),
		.io_dmem_req_ready                                  (io_dmem_req_ready                                  ),
		.io_dmem_req_valid                                  (io_dmem_req_valid                                  ),
		.io_dmem_resp_bits_data                             (io_dmem_resp_bits_data                             ),
		.io_dmem_resp_bits_data_word_bypass                 (io_dmem_resp_bits_data_word_bypass                 ),
		.io_dmem_resp_bits_has_data                         (io_dmem_resp_bits_has_data                         ),
		.io_dmem_resp_bits_replay                           (io_dmem_resp_bits_replay                           ),
		.io_dmem_resp_bits_tag                              (io_dmem_resp_bits_tag                              ),
		.io_dmem_resp_bits_typ                              (io_dmem_resp_bits_typ                              ),
		.io_dmem_resp_valid                                 (io_dmem_resp_valid                                 ),
		.io_dmem_s1_data_data                               (io_dmem_s1_data_data                               ),
		.io_dmem_s1_data_mask                               (io_dmem_s1_data_mask                               ),
		.io_dmem_s1_kill                                    (io_dmem_s1_kill                                    ),
		.io_dmem_s2_nack                                    (io_dmem_s2_nack                                    ),
		.io_dmem_s2_xcpt_ae_ld                              (io_dmem_s2_xcpt_ae_ld                              ),
		.io_dmem_s2_xcpt_ae_st                              (io_dmem_s2_xcpt_ae_st                              ),
		.io_dmem_s2_xcpt_ma_ld                              (io_dmem_s2_xcpt_ma_ld                              ),
		.io_dmem_s2_xcpt_ma_st                              (io_dmem_s2_xcpt_ma_st                              ),
		.io_dmem_s2_xcpt_pf_ld                              (io_dmem_s2_xcpt_pf_ld                              ),
		.io_dmem_s2_xcpt_pf_st                              (io_dmem_s2_xcpt_pf_st                              ),
		.io_fpu_dec_ren1                                    (io_fpu_dec_ren1                                    ),
		.io_fpu_dec_ren2                                    (io_fpu_dec_ren2                                    ),
		.io_fpu_dec_ren3                                    (io_fpu_dec_ren3                                    ),
		.io_fpu_dec_wen                                     (io_fpu_dec_wen                                     ),
		.io_fpu_dmem_resp_data                              (io_fpu_dmem_resp_data                              ),
		.io_fpu_dmem_resp_tag                               (io_fpu_dmem_resp_tag                               ),
		.io_fpu_dmem_resp_type                              (io_fpu_dmem_resp_type                              ),
		.io_fpu_dmem_resp_val                               (io_fpu_dmem_resp_val                               ),
		.io_fpu_fcsr_flags_bits                             (io_fpu_fcsr_flags_bits                             ),
		.io_fpu_fcsr_flags_valid                            (io_fpu_fcsr_flags_valid                            ),
		.io_fpu_fcsr_rdy                                    (io_fpu_fcsr_rdy                                    ),
		.io_fpu_fcsr_rm                                     (io_fpu_fcsr_rm                                     ),
		.io_fpu_fromint_data                                (io_fpu_fromint_data                                ),
		.io_fpu_illegal_rm                                  (io_fpu_illegal_rm                                  ),
		.io_fpu_inst                                        (io_fpu_inst                                        ),
		.io_fpu_killm                                       (io_fpu_killm                                       ),
		.io_fpu_killx                                       (io_fpu_killx                                       ),
		.io_fpu_nack_mem                                    (io_fpu_nack_mem                                    ),
		.io_fpu_sboard_clr                                  (io_fpu_sboard_clr                                  ),
		.io_fpu_sboard_clra                                 (io_fpu_sboard_clra                                 ),
		.io_fpu_sboard_set                                  (io_fpu_sboard_set                                  ),
		.io_fpu_store_data                                  (io_fpu_store_data                                  ),
		.io_fpu_toint_data                                  (io_fpu_toint_data                                  ),
		.io_fpu_valid                                       (io_fpu_valid                                       ),
		.io_hartid                                          (io_hartid                                          ),
		.io_imem_bht_update_bits_mispredict                 (io_imem_bht_update_bits_mispredict                 ),
		.io_imem_bht_update_bits_pc                         (io_imem_bht_update_bits_pc                         ),
		.io_imem_bht_update_bits_prediction_bits_bht_history(io_imem_bht_update_bits_prediction_bits_bht_history),
		.io_imem_bht_update_bits_prediction_bits_bht_value  (io_imem_bht_update_bits_prediction_bits_bht_value  ),
		.io_imem_bht_update_bits_prediction_valid           (io_imem_bht_update_bits_prediction_valid           ),
		.io_imem_bht_update_bits_taken                      (io_imem_bht_update_bits_taken                      ),
		.io_imem_bht_update_valid                           (io_imem_bht_update_valid                           ),
		.io_imem_btb_update_bits_br_pc                      (io_imem_btb_update_bits_br_pc                      ),
		.io_imem_btb_update_bits_cfiType                    (io_imem_btb_update_bits_cfiType                    ),
		.io_imem_btb_update_bits_isValid                    (io_imem_btb_update_bits_isValid                    ),
		.io_imem_btb_update_bits_pc                         (io_imem_btb_update_bits_pc                         ),
		.io_imem_btb_update_bits_prediction_bits_bht_history(io_imem_btb_update_bits_prediction_bits_bht_history),
		.io_imem_btb_update_bits_prediction_bits_bht_value  (io_imem_btb_update_bits_prediction_bits_bht_value  ),
		.io_imem_btb_update_bits_prediction_bits_entry      (io_imem_btb_update_bits_prediction_bits_entry      ),
		.io_imem_btb_update_bits_prediction_valid           (io_imem_btb_update_bits_prediction_valid           ),
		.io_imem_btb_update_valid                           (io_imem_btb_update_valid                           ),
		.io_imem_flush_icache                               (io_imem_flush_icache                               ),
		.io_imem_req_bits_pc                                (io_imem_req_bits_pc                                ),
		.io_imem_req_bits_speculative                       (io_imem_req_bits_speculative                       ),
		.io_imem_req_valid                                  (io_imem_req_valid                                  ),
		.io_imem_resp_bits_ae                               (io_imem_resp_bits_ae                               ),
		.io_imem_resp_bits_btb_bits_bht_history             (io_imem_resp_bits_btb_bits_bht_history             ),
		.io_imem_resp_bits_btb_bits_bht_value               (io_imem_resp_bits_btb_bits_bht_value               ),
		.io_imem_resp_bits_btb_bits_bridx                   (io_imem_resp_bits_btb_bits_bridx                   ),
		.io_imem_resp_bits_btb_bits_entry                   (io_imem_resp_bits_btb_bits_entry                   ),
		.io_imem_resp_bits_btb_bits_taken                   (io_imem_resp_bits_btb_bits_taken                   ),
		.io_imem_resp_bits_btb_valid                        (io_imem_resp_bits_btb_valid                        ),
		.io_imem_resp_bits_data                             (io_imem_resp_bits_data                             ),
		.io_imem_resp_bits_pc                               (io_imem_resp_bits_pc                               ),
		.io_imem_resp_bits_pf                               (io_imem_resp_bits_pf                               ),
		.io_imem_resp_bits_replay                           (io_imem_resp_bits_replay                           ),
		.io_imem_resp_ready                                 (io_imem_resp_ready                                 ),
		.io_imem_resp_valid                                 (io_imem_resp_valid                                 ),
		.io_imem_sfence_bits_rs1                            (io_imem_sfence_bits_rs1                            ),
		.io_imem_sfence_bits_rs2                            (io_imem_sfence_bits_rs2                            ),
		.io_imem_sfence_valid                               (io_imem_sfence_valid                               ),
		.io_interrupts_debug                                (io_interrupts_debug                                ),
		.io_interrupts_meip                                 (io_interrupts_meip                                 ),
		.io_interrupts_msip                                 (io_interrupts_msip                                 ),
		.io_interrupts_mtip                                 (io_interrupts_mtip                                 ),
		.io_interrupts_seip                                 (io_interrupts_seip                                 ),
		.io_ptw_invalidate                                  (io_ptw_invalidate                                  ),
		.io_ptw_pmp_0_addr                                  (io_ptw_pmp_0_addr                                  ),
		.io_ptw_pmp_0_cfg_a                                 (io_ptw_pmp_0_cfg_a                                 ),
		.io_ptw_pmp_0_cfg_l                                 (io_ptw_pmp_0_cfg_l                                 ),
		.io_ptw_pmp_0_cfg_r                                 (io_ptw_pmp_0_cfg_r                                 ),
		.io_ptw_pmp_0_cfg_w                                 (io_ptw_pmp_0_cfg_w                                 ),
		.io_ptw_pmp_0_cfg_x                                 (io_ptw_pmp_0_cfg_x                                 ),
		.io_ptw_pmp_0_mask                                  (io_ptw_pmp_0_mask                                  ),
		.io_ptw_pmp_1_addr                                  (io_ptw_pmp_1_addr                                  ),
		.io_ptw_pmp_1_cfg_a                                 (io_ptw_pmp_1_cfg_a                                 ),
		.io_ptw_pmp_1_cfg_l                                 (io_ptw_pmp_1_cfg_l                                 ),
		.io_ptw_pmp_1_cfg_r                                 (io_ptw_pmp_1_cfg_r                                 ),
		.io_ptw_pmp_1_cfg_w                                 (io_ptw_pmp_1_cfg_w                                 ),
		.io_ptw_pmp_1_cfg_x                                 (io_ptw_pmp_1_cfg_x                                 ),
		.io_ptw_pmp_1_mask                                  (io_ptw_pmp_1_mask                                  ),
		.io_ptw_pmp_2_addr                                  (io_ptw_pmp_2_addr                                  ),
		.io_ptw_pmp_2_cfg_a                                 (io_ptw_pmp_2_cfg_a                                 ),
		.io_ptw_pmp_2_cfg_l                                 (io_ptw_pmp_2_cfg_l                                 ),
		.io_ptw_pmp_2_cfg_r                                 (io_ptw_pmp_2_cfg_r                                 ),
		.io_ptw_pmp_2_cfg_w                                 (io_ptw_pmp_2_cfg_w                                 ),
		.io_ptw_pmp_2_cfg_x                                 (io_ptw_pmp_2_cfg_x                                 ),
		.io_ptw_pmp_2_mask                                  (io_ptw_pmp_2_mask                                  ),
		.io_ptw_pmp_3_addr                                  (io_ptw_pmp_3_addr                                  ),
		.io_ptw_pmp_3_cfg_a                                 (io_ptw_pmp_3_cfg_a                                 ),
		.io_ptw_pmp_3_cfg_l                                 (io_ptw_pmp_3_cfg_l                                 ),
		.io_ptw_pmp_3_cfg_r                                 (io_ptw_pmp_3_cfg_r                                 ),
		.io_ptw_pmp_3_cfg_w                                 (io_ptw_pmp_3_cfg_w                                 ),
		.io_ptw_pmp_3_cfg_x                                 (io_ptw_pmp_3_cfg_x                                 ),
		.io_ptw_pmp_3_mask                                  (io_ptw_pmp_3_mask                                  ),
		.io_ptw_pmp_4_addr                                  (io_ptw_pmp_4_addr                                  ),
		.io_ptw_pmp_4_cfg_a                                 (io_ptw_pmp_4_cfg_a                                 ),
		.io_ptw_pmp_4_cfg_l                                 (io_ptw_pmp_4_cfg_l                                 ),
		.io_ptw_pmp_4_cfg_r                                 (io_ptw_pmp_4_cfg_r                                 ),
		.io_ptw_pmp_4_cfg_w                                 (io_ptw_pmp_4_cfg_w                                 ),
		.io_ptw_pmp_4_cfg_x                                 (io_ptw_pmp_4_cfg_x                                 ),
		.io_ptw_pmp_4_mask                                  (io_ptw_pmp_4_mask                                  ),
		.io_ptw_pmp_5_addr                                  (io_ptw_pmp_5_addr                                  ),
		.io_ptw_pmp_5_cfg_a                                 (io_ptw_pmp_5_cfg_a                                 ),
		.io_ptw_pmp_5_cfg_l                                 (io_ptw_pmp_5_cfg_l                                 ),
		.io_ptw_pmp_5_cfg_r                                 (io_ptw_pmp_5_cfg_r                                 ),
		.io_ptw_pmp_5_cfg_w                                 (io_ptw_pmp_5_cfg_w                                 ),
		.io_ptw_pmp_5_cfg_x                                 (io_ptw_pmp_5_cfg_x                                 ),
		.io_ptw_pmp_5_mask                                  (io_ptw_pmp_5_mask                                  ),
		.io_ptw_pmp_6_addr                                  (io_ptw_pmp_6_addr                                  ),
		.io_ptw_pmp_6_cfg_a                                 (io_ptw_pmp_6_cfg_a                                 ),
		.io_ptw_pmp_6_cfg_l                                 (io_ptw_pmp_6_cfg_l                                 ),
		.io_ptw_pmp_6_cfg_r                                 (io_ptw_pmp_6_cfg_r                                 ),
		.io_ptw_pmp_6_cfg_w                                 (io_ptw_pmp_6_cfg_w                                 ),
		.io_ptw_pmp_6_cfg_x                                 (io_ptw_pmp_6_cfg_x                                 ),
		.io_ptw_pmp_6_mask                                  (io_ptw_pmp_6_mask                                  ),
		.io_ptw_pmp_7_addr                                  (io_ptw_pmp_7_addr                                  ),
		.io_ptw_pmp_7_cfg_a                                 (io_ptw_pmp_7_cfg_a                                 ),
		.io_ptw_pmp_7_cfg_l                                 (io_ptw_pmp_7_cfg_l                                 ),
		.io_ptw_pmp_7_cfg_r                                 (io_ptw_pmp_7_cfg_r                                 ),
		.io_ptw_pmp_7_cfg_w                                 (io_ptw_pmp_7_cfg_w                                 ),
		.io_ptw_pmp_7_cfg_x                                 (io_ptw_pmp_7_cfg_x                                 ),
		.io_ptw_pmp_7_mask                                  (io_ptw_pmp_7_mask                                  ),
		.io_ptw_ptbr_asid                                   (io_ptw_ptbr_asid                                   ),
		.io_ptw_ptbr_mode                                   (io_ptw_ptbr_mode                                   ),
		.io_ptw_ptbr_ppn                                    (io_ptw_ptbr_ppn                                    ),
		.io_ptw_status_dprv                                 (io_ptw_status_dprv                                 ),
		.io_ptw_status_mxr                                  (io_ptw_status_mxr                                  ),
		.io_ptw_status_prv                                  (io_ptw_status_prv                                  ),
		.io_ptw_status_sum                                  (io_ptw_status_sum                                  ),
		.io_rocc_cmd_ready                                  (io_rocc_cmd_ready                                  ),
		.io_rocc_cmd_valid                                  (io_rocc_cmd_valid                                  ),
		.io_rocc_interrupt                                  (io_rocc_interrupt                                  ),
		.reset                                              (reset                                              ),
		.rvfi_insn                                          (rvfi_insn                                          ),
		.rvfi_mem_addr                                      (rvfi_mem_addr                                      ),
		.rvfi_mem_rdata                                     (rvfi_mem_rdata                                     ),
		.rvfi_mem_rmask                                     (rvfi_mem_rmask                                     ),
		.rvfi_mem_wdata                                     (rvfi_mem_wdata                                     ),
		.rvfi_mem_wmask                                     (rvfi_mem_wmask                                     ),
		.rvfi_order                                         (rvfi_order                                         ),
		.rvfi_pc_rdata                                      (rvfi_pc_rdata                                      ),
		.rvfi_pc_wdata                                      (rvfi_pc_wdata                                      ),
		.rvfi_rd_addr                                       (rvfi_rd_addr                                       ),
		.rvfi_rd_wdata                                      (rvfi_rd_wdata                                      ),
		.rvfi_rs1_addr                                      (rvfi_rs1_addr                                      ),
		.rvfi_rs1_rdata                                     (rvfi_rs1_rdata                                     ),
		.rvfi_rs2_addr                                      (rvfi_rs2_addr                                      ),
		.rvfi_rs2_rdata                                     (rvfi_rs2_rdata                                     ),
		.rvfi_trap                                          (rvfi_trap                                          ),
		.rvfi_valid                                         (rvfi_valid                                         ),
	);
endmodule
